library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DDS_CTRL_v1_0 is
	generic (
		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH	: integer	:= 32;
		C_S00_AXI_ADDR_WIDTH	: integer	:= 6
	);
	port (
		-- Users to add ports here
		CUR_PROF        : in std_logic_vector(1023 downto 0);
		NXT_PROF        : in std_logic_vector(1023 downto 0);
        en_zond         : in std_logic;
        str_pn          : in std_logic;
        str_prd         : in std_logic;
        clk_dds         : in std_logic;
--        dds_io_upd_sinh : in std_logic;
        
        D               : out std_logic_vector(31 downto 0);
        F               : out std_logic_vector(3 downto 0);
        PS              : out std_logic_vector(2 downto 0);
        pwdwn           : out std_logic;
        rst             : out std_logic;
        osk_in          : in std_logic;
        osk_out         : out std_logic;
        drctrl_in       : in std_logic;
        drctrl_out      : out std_logic;
        drhold_in       : in std_logic;
        drhold_out      : out std_logic;
        drover_in       : in std_logic;
        drover_out      : out std_logic;
        io_upd_in       : in std_logic;
        io_upd_out      : out std_logic;
        sinc_out        : out std_logic;
        sinc_in         : in std_logic;
        dir             : out std_logic;

		-- User ports ends
		-- Do not modify the ports beyond this line


		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk	: in std_logic;
		s00_axi_aresetn	: in std_logic;
		s00_axi_awaddr	: in std_logic_vector(5 downto 0);
		s00_axi_awprot	: in std_logic_vector(2 downto 0);
		s00_axi_awvalid	: in std_logic;
		s00_axi_awready	: out std_logic;
		s00_axi_wdata	: in std_logic_vector(31 downto 0);
		s00_axi_wstrb	: in std_logic_vector(3 downto 0);
		s00_axi_wvalid	: in std_logic;
		s00_axi_wready	: out std_logic;
		s00_axi_bresp	: out std_logic_vector(1 downto 0);
		s00_axi_bvalid	: out std_logic;
		s00_axi_bready	: in std_logic;
		s00_axi_araddr	: in std_logic_vector(5 downto 0);
		s00_axi_arprot	: in std_logic_vector(2 downto 0);
		s00_axi_arvalid	: in std_logic;
		s00_axi_arready	: out std_logic;
		s00_axi_rdata	: out std_logic_vector(31 downto 0);
		s00_axi_rresp	: out std_logic_vector(1 downto 0);
		s00_axi_rvalid	: out std_logic;
		s00_axi_rready	: in std_logic
	);
end DDS_CTRL_v1_0;

architecture arch_imp of DDS_CTRL_v1_0 is

	-- component declaration
	component DDS_CTRL_v1_0_S00_AXI is
		port (		
		
		CUR_PROF        : in std_logic_vector(1023 downto 0);
		NXT_PROF        : in std_logic_vector(1023 downto 0);

        en_zond         : in std_logic;
        str_pn          : in std_logic;
        str_prd         : in std_logic;
        clk_dds         : in std_logic;
--        dds_io_upd_sinh : in std_logic;
        
        D               : out std_logic_vector(31 downto 0);
        F               : out std_logic_vector(3 downto 0);
        PS              : out std_logic_vector(2 downto 0);
        pwdwn           : out std_logic;
        rst             : out std_logic;
        osk_in          : in std_logic;
        osk_out         : out std_logic;
        drctrl_in       : in std_logic;
        drctrl_out      : out std_logic;
        drhold_in       : in std_logic;
        drhold_out      : out std_logic;
        drover_in       : in std_logic;
        drover_out      : out std_logic;
        io_upd_in       : in std_logic;
        io_upd_out      : out std_logic;
        sinc_out        : out std_logic;
        sinc_in         : in std_logic;
        dir             : out std_logic;

		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(5 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(31 downto 0);
		S_AXI_WSTRB	: in std_logic_vector(3 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(5 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(31 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component DDS_CTRL_v1_0_S00_AXI;

begin

-- Instantiation of Axi Bus Interface S00_AXI
DDS_CTRL_v1_0_S00_AXI_inst : DDS_CTRL_v1_0_S00_AXI
	port map (		
		CUR_PROF => CUR_PROF,
		NXT_PROF => NXT_PROF,
        en_zond => en_zond,
        str_pn => str_pn,
        str_prd => str_prd,
        clk_dds => clk_dds,
--        dds_io_upd_sinh => dds_io_upd_sinh,
        
        D => D,
        F => F,
        PS => PS,

        pwdwn => pwdwn,
        rst => rst,
        osk_in => osk_in,
        osk_out => osk_out,
        drctrl_in => drctrl_in,
        drctrl_out => drctrl_out,
        drhold_in => drhold_in,
        drhold_out => drhold_out,
        drover_in => drover_in,
        drover_out => drover_out,
        io_upd_in => io_upd_in,
        io_upd_out => io_upd_out,
        sinc_out => sinc_out,
        sinc_in => sinc_in,
        dir => dir,
		
		
		S_AXI_ACLK	=> s00_axi_aclk,
		S_AXI_ARESETN	=> s00_axi_aresetn,
		S_AXI_AWADDR	=> s00_axi_awaddr,
		S_AXI_AWPROT	=> s00_axi_awprot,
		S_AXI_AWVALID	=> s00_axi_awvalid,
		S_AXI_AWREADY	=> s00_axi_awready,
		S_AXI_WDATA	=> s00_axi_wdata,
		S_AXI_WSTRB	=> s00_axi_wstrb,
		S_AXI_WVALID	=> s00_axi_wvalid,
		S_AXI_WREADY	=> s00_axi_wready,
		S_AXI_BRESP	=> s00_axi_bresp,
		S_AXI_BVALID	=> s00_axi_bvalid,
		S_AXI_BREADY	=> s00_axi_bready,
		S_AXI_ARADDR	=> s00_axi_araddr,
		S_AXI_ARPROT	=> s00_axi_arprot,
		S_AXI_ARVALID	=> s00_axi_arvalid,
		S_AXI_ARREADY	=> s00_axi_arready,
		S_AXI_RDATA	=> s00_axi_rdata,
		S_AXI_RRESP	=> s00_axi_rresp,
		S_AXI_RVALID	=> s00_axi_rvalid,
		S_AXI_RREADY	=> s00_axi_rready
	);

	-- Add user logic here

	-- User logic ends

end arch_imp;
